`define SET_TIME_CMD      0

`define SET_ALARM_0_CMD   1
`define UNSET_ALARM_0_CMD 2

`define SET_ALARM_1_CMD   3
`define UNSET_ALARM_1_CMD 4

`define SET_ALARM_2_CMD   5
`define UNSET_ALARM_2_CMD 6

`define SET_ALARM_3_CMD   7
`define UNSET_ALARM_3_CMD 8

`define SET_ALARM_4_CMD   9
`define UNSET_ALARM_4_CMD 10

`define SET_ALARM_5_CMD   11
`define UNSET_ALARM_5_CMD 12

`define SET_ALARM_6_CMD   13
`define UNSET_ALARM_6_CMD 14

`define CMD_CNT 15
