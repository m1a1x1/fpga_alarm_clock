`define MONTH_CNT 12

`define JAN_DAYS_CNT 31
`define FEB_DAYS_CNT 28
`define FEB_LEAP_DAYS_CNT 29
`define MAR_DAYS_CNT 31
`define APR_DAYS_CNT 30
`define MAY_DAYS_CNT 31
`define JUNE_DAYS_CNT 30
`define JULY_DAYS_CNT 31
`define AUG_DAYS_CNT 31
`define SEPT_DAYS_CNT 30
`define OCT_DAYS_CNT 31
`define NOV_DAYS_CNT 30
`define DEC_DAYS_CNT 31     
