`define BLACK      3'b000
`define RED        3'b001
`define GREEN      3'b010
`define YELLOW     3'b011
`define BLUE       3'b100
`define PINK       3'b101
`define LIGHT_BLUE 3'b110
`define WIGHT      3'b111


